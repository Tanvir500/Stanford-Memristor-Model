`include "constants.vams"
`include "disciplines.vams"
module mem_stanford1(t,b);
    electrical t , b ;
    inout t , b ;

    parameter real a = 0.25e-9 ;       // unit: m  distance between adjacent oxygen vacancy 
    parameter real f = 1e13 ;          // unit: HZ  vibration frequency of oxygen atom in VO
    parameter real Ea = 0.7 ;          // unit: ev  average active energy of VO
    parameter real Eh = 1.12 ;          // unit: ev    hopping barrier of oxygen ion (O2-)     
    parameter real Ei = 0.82 ;          // unit: ev   energy barrier between the electrode and oxide
    parameter real r = 1.5 ;           // enhancement factor of external voltage
    parameter real alphah = 0.75e-9 ;  // unit: m   enhancement factor in lower Ea & Eh
    parameter real alpha = 0.75e-9 ;   // unit: m    enhancement factor in lower Ea & Eh
    parameter real Z = 1 ;
    parameter real XT = 0.4e-9 ;       // unit: m          
    parameter real VT = 0.4 ;          // unit: V
    parameter real L0 = 3e-9 ;         // unit: m     L0 is defined as the initial fixed length of the RRAM switching layer
    parameter real x0 = 3e-9 ;         // unit: m    x0 is defined as the initial length of gap region during both SET/RESET (for SET: x0=L0)
    parameter real w0 = 0.5e-9 ;       // unit: m    initial CF width
    parameter real WCF = 5e-9 ;        // unit: m   fixed width of the RRAM switching layer
    parameter real weff = 0.5e-9 ;     // unit: m     effective CF extending width
    parameter real I0 = 1e13 ;         // unit: A/m^2    hopping current density in the gap region
    parameter real rou = 1.9635e-5 ;   // unit: ohm*m   resistivity of the formed conductive filament (CF)
    parameter real pi = 3.1415926 ;    
    parameter real Rth = 5e5 ;         // unit: K/W   effective thermal resistance
    parameter real Kb = 8.61733e-5 ;   // unit: ev/K
    parameter real T0 = 300 ;          // unit: K   ambient temperature
    parameter real switch = 1  ;          // switch = 1: variation-included ; switch = 0: no variations
    parameter real deltaGap = 4e-5 ;     // gap distance variation amplitude
    parameter real deltaCF     = 1e-4 ;  // filament radius variation amplitude
    parameter real crit_x = 0.5e-9 ;     // decided by measured variation amplitude
    parameter real user_seed = 0 ;       // specified user seed for random number generator 
    
    real Temp=T0 ;
    real dxr1 ;
    real dxr2 ;
    real dxs ;
    real dx=0 ;   
    real dw=0 ;
    real x=x0 ;    
    real w=w0 ;
    real RCF ;
    real Vg ;
    real I1 ;

    integer rand_seed_set  ;
    integer rand_seed_reset ;
    real cf_random_ddt ;       
    real gap_random_ddt ;

    analog 
    begin
        Temp = T0 + abs(I(t,b) * V(t,b)) * Rth ;
        I1 = I0*pi*(WCF*WCF/4-w*w/4)*exp(-L0/XT)*sinh(V(t,b)/VT) ;
        RCF = rou*(L0-x)/(pi*w*w/4) ;            
        Vg = V(t,b) - (I(t,b)-I1)*RCF ;

        if ( V(t,b) > 0 ) 
        begin
            if ( x > 0 )
            begin
                dxs = -a*f*exp(-(Ea-Vg*alpha*Z/x)/(Kb*Temp)) ;
                if ( abs(dxs) <= 1e2 )
                begin
                    dx = dxs ;
                end
                else
                begin
                    dx = -1e2 ;
                end
            end
            else if ( x <= 0 )
            begin
                dx = 0 ;           
            end
            
            if ( w < WCF )
            begin
                dw = (x>0)*0 + (x<=0)*(weff+pow(weff,2)/(2*w))*f*exp(-(Ea-V(t,b)*alpha*Z/L0)/(Kb*Temp)) ;
                if ( dw > 1e2 )
                begin   
                    dw = 1e2 ;
                end
            end
            else if ( w >= WCF)
                dw = 0 ;
                
        end
        else if ( V(t,b) < 0 )
        begin
            dw = 0 ;
            if ( x <= 0 )   
            begin
                dxr1 = a*f*exp(-(Ei+r*Z*Vg)/(Kb*Temp)) ;
                dx = dxr1 ;
            end
            else if ( x > 0 )
            begin
                if ( x < L0 )
                begin
                    dxr1 = a*f*exp(-(Ei+r*Z*Vg)/(Kb*Temp)) ;
                    dxr2 = a*f*exp(-Eh/(Kb*Temp))*sinh(alphah*Z*-1*Vg/(x*Kb*Temp)) ;
                    dx = (dxr1<dxr2)*dxr1 + (dxr2<=dxr1)*dxr2 ;
                end
                else if ( x >= L0 )  
                begin
                    dx = 0 ;
                end                 
            end 
        end
        else if ( V(t,b) == 0 )
        begin
            dx = 0 ;
            dw = 0 ;
        end
    
        if ( V(t,b) == 0 )
        begin
            I(t,b) <+ 0 ;
        end
        else if ( V(t,b) > 0 )
        begin
            if ( x > 0 )
            begin
                I(t,b) <+ I1 + I0*pi*(w*w/4)*exp(-x/XT)*sinh(Vg/VT) ;
            end
            else if ( x <= 0 )
            begin
                I(t,b) <+ I1 + V(t,b)/(rou*L0/(pi*w*w/4)) ;   
            end
        end
        else if ( V(t,b) < 0 )
        begin
            I(t,b) <+ I1 + I0*pi*(w*w/4)*exp(-x/XT)*sinh(Vg/VT) ;
        end

        if ( switch == 1 )
        begin   
            if ( V(t,b) > 0 )
            begin
                if ( dw == 0 )
                begin
                    cf_random_ddt = 0 ;
                end
                else
                begin
                    rand_seed_set = $random + user_seed ;
                    cf_random_ddt = $rdist_normal(rand_seed_set,0,1) * deltaCF ;
                end
            end
            else if ( V(t,b) < 0 )
            begin
                if ( x < crit_x )
                begin
                    gap_random_ddt = 0 ;
                end
                else if ( x >= crit_x )
                begin
                    rand_seed_reset = $random + user_seed ;
                    gap_random_ddt = $rdist_normal(rand_seed_reset,0,1) * deltaGap ;
                end
            end
            else
            begin
                gap_random_ddt = 0 ;
                cf_random_ddt = 0 ;
            end
        end
        else
        begin
            gap_random_ddt = 0 ;
            cf_random_ddt = 0 ;
        end
        
        x = idt(dx+gap_random_ddt,x0) ;
        w = idt(dw+cf_random_ddt,w0) ;
    
        if ( x < 0 ) 
        begin
            x = 0 ;
        end
        if ( x > L0 )
        begin
            x = L0 ;
        end
        
        if ( w > WCF ) 
        begin
            w = WCF ;
        end
    end

endmodule


